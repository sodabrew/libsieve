require ["reject"];
reject text:
I don't like your face
Or your dog.
   Or anything else.
..
.
;
