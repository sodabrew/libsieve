require "vacation";

vacation :days 2 
      :subject "I'm just not here"
      "Look folks, I'm not here. Period. Go away!";

