discard;
