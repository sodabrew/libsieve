require ["fileinto"];
asdf
asdf
asdf
asdf
asdf
;
