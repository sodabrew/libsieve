require "vacation";

vacation :subject "I'm just not here" 
:days 2
 :handle "foo12345"
	:from "vacation@localhost"
"Look folks, I'm not here. Period. Go away!";

