
if header :contains "Subject" "$${hex:24 24}" {
	discard;
}

