require ["fileinto", "reject"];

fileinto "Rejected Messages";

reject "I don't like you.";
